//======================================================================================= 
// TITLE : Result receiver for Sharp LR35902 ALU
// DESCRIPTION : 
// 
// Read result from the Sharp LR35902 ALU each clock cycle and send result packet to scoreboard
//
// FILE : Monitor.sv
//======================================================================================= 
// CREATION 
// DATE AUTHOR PROJECT REVISION 
// 2015/07/28 Etienne Gauthier 
//======================================================================================= 
// MODIFICATION HISTORY 
// DATE AUTHOR PROJECT REVISION COMMENTS 
// 2018/01/21 Etienne Gauthier Ajout du format du module moniteur
//======================================================================================= 
`include "Sharp_LR35902_alu_opcodes.v"

module Monitor (Interface_to_alu intf_dut);

	// ### À compléter ###

endmodule